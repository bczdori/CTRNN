** Profile: "teljes_aramkor-telj_aramkor3"  [ C:\Users\Public\babdo\orcad_projects\article_circuit3\article_circuit3-pspicefiles\teljes_aramkor\telj_aramkor3.sim ] 

** Creating circuit file "telj_aramkor3.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
* From [PSPICE NETLIST] section of C:\SPB_Data\cdssetup\OrCAD_PSpice/16.6.0/PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 5m 0 500n SKIPBP 
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\teljes_aramkor.net" 


.END
